library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity av_master_simple_tb is
	end entity av_master_simple_tb;
	
architecture bench of av_master_simple_tb is
begin 
	end architecture bench;