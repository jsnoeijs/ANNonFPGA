library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


entity gru_ppl_tb is
	end entity gru_ppl_tb;
	
architecture bench of gru_ppl_tb is
begin 
	end architecture bench;