library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity activation is
	end entity activation;
	
architecture simple of activation is
begin
	end architecture simple;