library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity av_slave is
	end entity av_slave;
	
architecture simple of av_slave is
begin
	end architecture simple;
