library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity av_master is
	end entity av_master;
	
architecture simple of av_master is
begin
	end architecture simple;
